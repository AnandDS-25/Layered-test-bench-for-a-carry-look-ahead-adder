interface intf();
  
  logic [31:0]a;
  logic [31:0]b;
  logic cin;
  logic [31:0]s;
  logic cout;
  
endinterface