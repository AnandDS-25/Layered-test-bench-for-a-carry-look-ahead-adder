module prop(input logic a,b, output logic p);
assign p=a|b;
endmodule